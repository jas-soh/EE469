// todo, create pipelined cpu
module Pipelined_CPU(reset, clk);
	input logic clk, reset;
endmodule


// This module is the execution stage.
// Controls passed on: MemWE, Mem2Reg, and RegWE.
module EX ();

endmodule
module ID_EX_reg ();

    // alu alu_operation (.A(Da), .B(ALUSrc_out), .cntrl(ALUOp), .result(ALU_out),
    //     negative(negFlag), .zero(ALUzeroFlag), .overflow(ovFlag), .carry_out_flag(cOutFlag));

    //input logic 

endmodule